version https://git-lfs.github.com/spec/v1
oid sha256:8dd989ca74750695d39095182c48a69eef555a2996d0c97ee2a0db9479cfd1d5
size 6430
