version https://git-lfs.github.com/spec/v1
oid sha256:b848390b6594fcc8d2eae6ab5e2a2e7bdc6c1d8d35ccd013b575c549139d4b06
size 1270
