version https://git-lfs.github.com/spec/v1
oid sha256:36857ff2b8bc3b681350eedd88a52e98b010c75d6718d3496eddce4951520d3b
size 1401
