version https://git-lfs.github.com/spec/v1
oid sha256:0248a9a08f0be4ef509ee234d4cc30f64afd14ff2838fd2179d147ed687c7bd8
size 2697
