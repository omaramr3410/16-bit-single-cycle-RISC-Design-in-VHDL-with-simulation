version https://git-lfs.github.com/spec/v1
oid sha256:1deccef29e4980a1ac7e3805b67b71b5bfbe6b1e5f3186fd26485e8dff57f46b
size 2484
