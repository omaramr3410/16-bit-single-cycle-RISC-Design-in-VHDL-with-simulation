version https://git-lfs.github.com/spec/v1
oid sha256:c640c9ce725c22dea4bafb0ebb764c4e2aa9895eac2a93720d8be566f0b2efb8
size 2717
