version https://git-lfs.github.com/spec/v1
oid sha256:259b7205d88c4b27e2f99ab2af974e352d7a38672cbe23e264d5b6101533ec2b
size 3250
