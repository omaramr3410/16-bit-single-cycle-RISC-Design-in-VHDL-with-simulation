version https://git-lfs.github.com/spec/v1
oid sha256:d65fd432ed8886b38e77e9e04c045ac37390f4496c16778eff7b1e3d359a175d
size 8054
