version https://git-lfs.github.com/spec/v1
oid sha256:e06e4df780e7f36fd28f494dfda907dd59bdae80a8e47b4b6330006c2abe5a79
size 3482
