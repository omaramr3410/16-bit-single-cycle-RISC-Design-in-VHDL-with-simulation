version https://git-lfs.github.com/spec/v1
oid sha256:072ee611872c97aba1bdb485d0dc5df76d525fb143783f47b820e6a830ae7958
size 2031
