version https://git-lfs.github.com/spec/v1
oid sha256:53bacd8cd1d883aa90ecb31e748e39f689a90787ae71ab88fbba58297f571f4f
size 1784
