version https://git-lfs.github.com/spec/v1
oid sha256:55974cfd1266209909fd3ecc4d8291964ebc8cd70acd44ee8b7c21759a0e0aea
size 1903
