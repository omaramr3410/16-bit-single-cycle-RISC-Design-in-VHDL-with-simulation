version https://git-lfs.github.com/spec/v1
oid sha256:053b1d9d2a1de40e146075f240fd93b39347467269accc66493cd276fb94c640
size 1892
