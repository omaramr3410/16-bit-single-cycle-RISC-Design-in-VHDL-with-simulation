version https://git-lfs.github.com/spec/v1
oid sha256:f4381a4653fd485c0621cf885622300e6ea592cade2fa08f13a5418893a3c7e5
size 3279
