version https://git-lfs.github.com/spec/v1
oid sha256:a0aa376391cf75fc293aeceb712c5eb012c013b3542b2922fc992f85d9b58d5c
size 2139
