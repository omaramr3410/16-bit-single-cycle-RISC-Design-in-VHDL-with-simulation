version https://git-lfs.github.com/spec/v1
oid sha256:8ca253e495b4b628c5dfdc0e1d21eabe2a64731ee281226f717d2ca0187ea06c
size 1906
