version https://git-lfs.github.com/spec/v1
oid sha256:4b928fec9b34f60829b8456f4873901020459e0f68cff04fea1be5c8965253eb
size 2599
