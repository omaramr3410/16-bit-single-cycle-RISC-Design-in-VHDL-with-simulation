version https://git-lfs.github.com/spec/v1
oid sha256:2e8763e41de69a6d71fde834cbaa16e19a9106cdd7b49e958276175267219563
size 5522
