version https://git-lfs.github.com/spec/v1
oid sha256:60ca2fe5c7a158a0095dc5889f2fa7ccfd8538f5fba57a77700d783036959297
size 6150
