version https://git-lfs.github.com/spec/v1
oid sha256:321679e61fadd211277c7ae23c246f27e2efbf5e6e444e72ee45bb1a0025c0d9
size 3245
