version https://git-lfs.github.com/spec/v1
oid sha256:256a4a2f48828aa688cfbf546d98097c18e9842a82269d1f36398cc996783c65
size 709
