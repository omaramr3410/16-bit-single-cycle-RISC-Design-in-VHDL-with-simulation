version https://git-lfs.github.com/spec/v1
oid sha256:5fcd8763b94b91086de6f93bb023f2dee0caf7803bd2c3d977ff35206b6a77f1
size 2628
