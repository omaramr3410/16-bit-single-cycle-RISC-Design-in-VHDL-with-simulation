version https://git-lfs.github.com/spec/v1
oid sha256:52597ee906047f3a6c7f3b3a0409f96b77d56afe9eda35300a91d99cd9dc1c47
size 1217
