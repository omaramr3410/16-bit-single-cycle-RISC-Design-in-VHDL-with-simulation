version https://git-lfs.github.com/spec/v1
oid sha256:f29b6a07cd4b828ca1ecea20249e542d94f3fde6fd598c1eaf4a826efb07d567
size 5747
