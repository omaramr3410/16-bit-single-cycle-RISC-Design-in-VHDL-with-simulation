version https://git-lfs.github.com/spec/v1
oid sha256:baa13ef89d59279fd62a6587c0603cada930f92da57a47c88abf91effb5492a4
size 6047
