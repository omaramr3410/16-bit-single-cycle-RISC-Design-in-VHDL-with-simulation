version https://git-lfs.github.com/spec/v1
oid sha256:57936bd7c913ee95fcf03859b550084562de5eb960b5f19c6e4739d04eb8f9d3
size 5555
