version https://git-lfs.github.com/spec/v1
oid sha256:01c05132180bea4b35df0405ab94b8e45047421b0d126a35ccf2aedfaec5f469
size 2191
