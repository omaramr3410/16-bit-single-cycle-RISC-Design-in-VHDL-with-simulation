version https://git-lfs.github.com/spec/v1
oid sha256:eaba2bc4916d30827189429bba698f58728a5040c0e34b2fd14599fd60ec5645
size 1426
