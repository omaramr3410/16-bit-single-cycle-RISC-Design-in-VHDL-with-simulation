version https://git-lfs.github.com/spec/v1
oid sha256:77fd99bd9c804219ab0ae8c4be1fbdb06ef9e664e710cf4e14ab35a7273b485d
size 6256
