version https://git-lfs.github.com/spec/v1
oid sha256:06d29989a005730a5fa933eadecc9d620e06d6d53419fc09c9ee3947c0fe2225
size 717
