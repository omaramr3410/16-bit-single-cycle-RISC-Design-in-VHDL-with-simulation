version https://git-lfs.github.com/spec/v1
oid sha256:ac13e6b4857773b5315a47e03b17b9dbf6617f05e00adadfa73105bbc60dc45f
size 2764
