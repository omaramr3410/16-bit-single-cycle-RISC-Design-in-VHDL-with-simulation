version https://git-lfs.github.com/spec/v1
oid sha256:0e3e99c5fbc1fde7b7a7672cd7fa8c59327247f1b8e428153ff028efc9c5d0d2
size 2424
