version https://git-lfs.github.com/spec/v1
oid sha256:d7d045716617f347b45f34b432e1038c2e1b9c2f2dc3fd7f424ed528a7aceea2
size 7043
