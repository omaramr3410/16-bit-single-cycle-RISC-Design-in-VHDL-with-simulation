version https://git-lfs.github.com/spec/v1
oid sha256:0b80e418c8cc97111c1d2f7f6394c5133b9415c17188adaf00d1b47f59646dc6
size 2507
