version https://git-lfs.github.com/spec/v1
oid sha256:e680ac46b2e48a58eff9e7bd9f5aea86bca56e8316f85df194cfa2d7c14b4e56
size 1247
