version https://git-lfs.github.com/spec/v1
oid sha256:492d0703848905f91eefe7fac4b1c10253dcff3700908488fb6f5e5476090fa7
size 393
