version https://git-lfs.github.com/spec/v1
oid sha256:fdd8304621d9ba89548b1cc2e4ba043d3fa658f42e1b936705c082aaa7397012
size 414
