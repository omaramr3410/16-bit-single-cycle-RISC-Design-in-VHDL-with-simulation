version https://git-lfs.github.com/spec/v1
oid sha256:185bbd4e6860ebef442fb60911ccbac82b0121fa3b5459085d9c65b0f4639983
size 2185
