version https://git-lfs.github.com/spec/v1
oid sha256:c61307c9a99de000660f6efb010b2d398338dfb3bd922fc3d2b0da3854784730
size 2217
