version https://git-lfs.github.com/spec/v1
oid sha256:7d420c854386864ee8077d71c6d54ca2fa11c412a4186d4968c03b990b2ef214
size 6631
