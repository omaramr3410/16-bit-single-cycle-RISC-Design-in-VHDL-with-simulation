version https://git-lfs.github.com/spec/v1
oid sha256:676f51cf7df0a630094e2abc2ce378db74011204a3cb49eab636f8bb4c30b1ef
size 1497
