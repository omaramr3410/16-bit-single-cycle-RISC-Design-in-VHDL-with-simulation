version https://git-lfs.github.com/spec/v1
oid sha256:671a5ab19885fa3b2ab52dfe7964ef926048cf1446ba5c53e0f143598a455ac7
size 2484
