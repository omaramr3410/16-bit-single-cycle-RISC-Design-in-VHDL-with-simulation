version https://git-lfs.github.com/spec/v1
oid sha256:9f51962645b80acfac2479822bfcf678f40af8e7469717ac63ce6a6532ffd9b6
size 682
