version https://git-lfs.github.com/spec/v1
oid sha256:9baa532b5faecf8c435c7038443a4428bc204f0bbd9ac80aaffa23dac2891590
size 1844
