version https://git-lfs.github.com/spec/v1
oid sha256:060a66ff1b4b2661cb0680d3439f4e95ce8d0d8b323e5e9b583ded5618e2b145
size 6155
