version https://git-lfs.github.com/spec/v1
oid sha256:24e1bfdc80160d8dc3da342bea4a8073b7bbc2b4cc5343228e4cb2a2e577ef81
size 1241
