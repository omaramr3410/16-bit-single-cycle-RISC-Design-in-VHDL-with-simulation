version https://git-lfs.github.com/spec/v1
oid sha256:28e18757053c1f9d6a78aa6fb53c654b8d3a244d90c76bdfc03ff4f91ce68d83
size 8107
