version https://git-lfs.github.com/spec/v1
oid sha256:fab05c922479502afd9f026b458b639af3f6c08d5cbabd86046bb9f29e6d1836
size 694
