version https://git-lfs.github.com/spec/v1
oid sha256:8a8a94cad50e637c238e4365d623c361395e6cc7ef64f8e31afda064bb46b2af
size 6051
