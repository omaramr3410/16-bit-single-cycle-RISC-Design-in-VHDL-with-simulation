version https://git-lfs.github.com/spec/v1
oid sha256:a3fd6d1e3e10674ddec5393c8b9a219ce36de1786f12dcf58a063ab73ec80496
size 7709
