version https://git-lfs.github.com/spec/v1
oid sha256:438b7547d794d5c20405399d64af708c688c38695cfee3c00688b0f555036c66
size 731
