version https://git-lfs.github.com/spec/v1
oid sha256:99477c94da756255c4eb8826503b657d5ba4d648b208347edc27121290f3c295
size 1087
