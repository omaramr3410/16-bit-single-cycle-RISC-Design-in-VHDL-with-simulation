version https://git-lfs.github.com/spec/v1
oid sha256:a77056d72b22e33977f8e61890574290cce1324ec4ac2319a2cdc9d32be8d033
size 3428
