version https://git-lfs.github.com/spec/v1
oid sha256:2c67c5f517df1363be2d7faa80a40db211a695b954c532534c305a3e69346b8f
size 1229
