version https://git-lfs.github.com/spec/v1
oid sha256:67d408fadb13988371e07306e7af9149f6ba8d7c853649d61e05bd78b67086ad
size 1827
