version https://git-lfs.github.com/spec/v1
oid sha256:2e9ee7a335882f1c2a576e96b50b0534b5b21a9fcdac2f7c581ab75ba9400f35
size 1988
