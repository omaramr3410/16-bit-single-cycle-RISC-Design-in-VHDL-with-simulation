version https://git-lfs.github.com/spec/v1
oid sha256:8fdb314c68511b846800a97a3eb0af9bd1f7a0bac18a4bd7835a350c0ca803c1
size 3443
