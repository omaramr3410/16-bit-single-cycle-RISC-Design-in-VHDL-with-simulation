version https://git-lfs.github.com/spec/v1
oid sha256:f3341eca8efd94411fea4e145ce8ead27a837b6fde92afddfd1989597a05ffdd
size 411
