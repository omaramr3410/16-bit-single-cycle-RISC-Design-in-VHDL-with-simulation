version https://git-lfs.github.com/spec/v1
oid sha256:762b99d4f5fb133108217b2251e3562a46f1590fcf304babad2e15cccd2ac7c9
size 2499
