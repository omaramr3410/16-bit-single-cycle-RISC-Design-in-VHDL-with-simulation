version https://git-lfs.github.com/spec/v1
oid sha256:bd3890736d8820cef39d803bd9c7a82126cd2d148336629098d1b15783ddd92c
size 2296
