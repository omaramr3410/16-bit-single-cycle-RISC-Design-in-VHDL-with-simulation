version https://git-lfs.github.com/spec/v1
oid sha256:3ae968b13dae3e3128085184ee28f89690a54af894d16ac96bf57c022ce92bb1
size 8219
