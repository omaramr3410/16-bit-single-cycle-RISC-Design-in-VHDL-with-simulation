version https://git-lfs.github.com/spec/v1
oid sha256:beb3a58d6b818d43219979d2c6cec8b86769774d939db1357f0ca5abbb726cf3
size 1422
