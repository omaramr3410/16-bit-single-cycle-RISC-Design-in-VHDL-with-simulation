version https://git-lfs.github.com/spec/v1
oid sha256:ae274643c281642c15826ba19f2ef553d7313427d35fc5e996a3832998a08ac3
size 1931
