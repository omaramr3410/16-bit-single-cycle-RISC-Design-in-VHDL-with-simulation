version https://git-lfs.github.com/spec/v1
oid sha256:653b6c39c5a5a4b6aabca0016884438924e1375fabb3095485b9f47f00859574
size 4827
