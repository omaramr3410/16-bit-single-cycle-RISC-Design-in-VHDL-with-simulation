version https://git-lfs.github.com/spec/v1
oid sha256:c41d8b9ee8e0a5f85ab652cc2e9f5a43233baf1d3f4cf217f7b54b87983d0b09
size 2151
