version https://git-lfs.github.com/spec/v1
oid sha256:1ffbab73acd361f9426420c399e5f4fa44df15e52b11cd466faf497d88e62b96
size 2564
