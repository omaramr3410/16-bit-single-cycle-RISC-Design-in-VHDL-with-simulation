version https://git-lfs.github.com/spec/v1
oid sha256:3c76daa759b5cbcc4dbfb1487933214e408249ed3d95100a808b1b259ef8be48
size 1240
