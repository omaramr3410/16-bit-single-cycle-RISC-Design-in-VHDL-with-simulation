version https://git-lfs.github.com/spec/v1
oid sha256:1c0f2c978cbbd3ba3b1ec63e786eccddc145ac50399f2669d200a9bdd16d6328
size 640
