version https://git-lfs.github.com/spec/v1
oid sha256:c053da91bc77d29a35ceb6d2d51fa63e1ab91de1f3bec8eb52757229d1e4b392
size 703
