version https://git-lfs.github.com/spec/v1
oid sha256:b7748cd8f6e9adc9fe205b9b6b7e87e664d4502192b8f28edf362aeb9478f3c5
size 2699
