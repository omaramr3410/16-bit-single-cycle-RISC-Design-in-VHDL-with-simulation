version https://git-lfs.github.com/spec/v1
oid sha256:9ddc89720796ee682f5ec1c59d16c9ad095c696ca412081584d8bb8445a7d2ed
size 8594
