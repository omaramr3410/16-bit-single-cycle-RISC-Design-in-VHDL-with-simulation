version https://git-lfs.github.com/spec/v1
oid sha256:c84b0dc3b7c959429f2582cf3e7b6ee05ac552b59d18dbe43a327566c3f7d077
size 7233
