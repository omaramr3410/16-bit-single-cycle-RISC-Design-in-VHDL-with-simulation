version https://git-lfs.github.com/spec/v1
oid sha256:d2e4ffeb548b890f776c8e16683797de25e35741e109f9c0400089ee250bd23e
size 1714
