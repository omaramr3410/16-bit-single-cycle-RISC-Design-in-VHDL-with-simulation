version https://git-lfs.github.com/spec/v1
oid sha256:8745ae3dae48b147a183205968f5b26bdc3f8be59548b5f768abfb004d932675
size 1284
