version https://git-lfs.github.com/spec/v1
oid sha256:da37f428fee89f8f9ca39a503d91b09354a12cd7778161734a720541169e389f
size 6991
