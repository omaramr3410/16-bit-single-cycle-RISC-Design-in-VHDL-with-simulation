version https://git-lfs.github.com/spec/v1
oid sha256:d00109a21b491569a12a3a613fc31d5642a027e5f457e2afd5b6c0f84e6fcb05
size 7046
