version https://git-lfs.github.com/spec/v1
oid sha256:5a170bb6033d22ca2b14c2f4849274fc09e7a0273c334a675d8f2658daa2703d
size 6943
