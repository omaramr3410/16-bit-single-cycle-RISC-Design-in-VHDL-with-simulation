version https://git-lfs.github.com/spec/v1
oid sha256:a9f9121ac56f8f2381f224e0cfd1e824ad51a7191c0591da203c67fa28faac9a
size 7131
