version https://git-lfs.github.com/spec/v1
oid sha256:2559a7c4094ea7a6eccc2107029cf1335e514afd1cec812430e663e5345ca92c
size 7271
