version https://git-lfs.github.com/spec/v1
oid sha256:e3670f7c0db13668515b41241386d6ed5975405bb367f16143f2c1622f3eb790
size 2399
