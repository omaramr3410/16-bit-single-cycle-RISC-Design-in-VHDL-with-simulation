version https://git-lfs.github.com/spec/v1
oid sha256:3e8e589c74734ccb4b4c0ad128b0a569f9d6c684ad080a132491d91a87bb7398
size 703
