version https://git-lfs.github.com/spec/v1
oid sha256:631dece8c019eb15eed8306aaa741b3d40f74f4be598ed4b55dbcdacb67c2d7d
size 5170
