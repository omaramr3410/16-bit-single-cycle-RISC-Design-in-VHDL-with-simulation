version https://git-lfs.github.com/spec/v1
oid sha256:1544b4d012e2d0f301147c0286adf15f7b72f41356f15a47e35de5f885abe37d
size 592
