version https://git-lfs.github.com/spec/v1
oid sha256:05cb39675bb1688e7d9ad1b2614b20da00ea90ec40c0cbd484c4eb5275e71c37
size 7041
