version https://git-lfs.github.com/spec/v1
oid sha256:e0adbe861428860cd2eff3a679d5c40c818f23bda583d7c01567e09b92487c20
size 5426
