version https://git-lfs.github.com/spec/v1
oid sha256:ca6702331ff0e4db8a6ea090bf6291a4f45578a1f466bd7eee02e891ab890519
size 3466
