version https://git-lfs.github.com/spec/v1
oid sha256:3f0c1a8491f0d62814db7da9405150130171722d95b7d5a6999cf0670c3d913b
size 1805
