version https://git-lfs.github.com/spec/v1
oid sha256:c86bb396c2df88d8f5c77619e0b8c06582c25792beb166082189972ac23392df
size 1763
