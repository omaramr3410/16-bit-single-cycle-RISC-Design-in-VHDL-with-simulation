version https://git-lfs.github.com/spec/v1
oid sha256:45af84927cda67d5b5798f9dca65c066db8aff8f42cd41e6ef121c46701afc83
size 1974
