version https://git-lfs.github.com/spec/v1
oid sha256:14cd02ae59154a38eb3978fbf2be2ef13589c31b2db9742f7000f1303e48a78d
size 5523
