version https://git-lfs.github.com/spec/v1
oid sha256:39e6f18e3e9f33464f1f369faefd99f6aae148fa8549b2bba92c88e0a9d107db
size 2030
