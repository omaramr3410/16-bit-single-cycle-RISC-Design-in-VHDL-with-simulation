version https://git-lfs.github.com/spec/v1
oid sha256:e606be83b8d212816d986a7715238ba3a34ba5987bc31e9b41431c508699518a
size 6429
