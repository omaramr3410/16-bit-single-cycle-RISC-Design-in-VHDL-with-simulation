version https://git-lfs.github.com/spec/v1
oid sha256:d9eff31f222bb5ab94888e7ab9e85bed0b41176a3eb4a96247d7b3a41e9f8b68
size 596
