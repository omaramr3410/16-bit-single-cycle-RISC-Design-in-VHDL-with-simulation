version https://git-lfs.github.com/spec/v1
oid sha256:0f489ebea09b7064e95c79140fdd79d0fa638699f1faf5d7616ae136a2a34426
size 1922
