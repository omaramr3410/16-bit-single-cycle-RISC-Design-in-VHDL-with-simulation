version https://git-lfs.github.com/spec/v1
oid sha256:29f0803c77c63c979fe1b6b2061bd2c35039e8d558124d0c520b64e29aa83602
size 3459
