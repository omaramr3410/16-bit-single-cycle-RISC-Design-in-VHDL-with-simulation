version https://git-lfs.github.com/spec/v1
oid sha256:a7c66b54367532e17b0c8fa0a9b2f541afa69e2cf5d975509af9534f47e6a1e9
size 9179
