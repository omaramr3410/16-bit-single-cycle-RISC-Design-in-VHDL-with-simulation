version https://git-lfs.github.com/spec/v1
oid sha256:5dbfb2a31f33a0dd8821dadae879e3f7292c27d019fe2009ce9b102c7e65ec26
size 1244
