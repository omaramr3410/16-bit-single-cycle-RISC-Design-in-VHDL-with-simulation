version https://git-lfs.github.com/spec/v1
oid sha256:1f63c6cc99a5c81f7809ba656757e93abf703eaf2354d2d2656ce24327872a81
size 2736
