version https://git-lfs.github.com/spec/v1
oid sha256:4fc6fd855e83e11934a8e03fb1f069548aaea25c7dc613b9fa1dffbaebde11a2
size 5630
