version https://git-lfs.github.com/spec/v1
oid sha256:628bc1498f570237e09b20c81fd350312a423f124af197cccc07dc58a65f08f0
size 1223
