version https://git-lfs.github.com/spec/v1
oid sha256:2447fc5248d5ddccb86519456af61b3da87f19da45f6e59b805615129031c897
size 668
