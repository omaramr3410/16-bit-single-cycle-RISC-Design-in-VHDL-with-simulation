version https://git-lfs.github.com/spec/v1
oid sha256:3d02add8d0dd4d44dc23272ff6358363a08874f7165c0c380d1c7399c634499e
size 2972
