version https://git-lfs.github.com/spec/v1
oid sha256:17633fee691e44fcb6787c1d9193186598e694d6644c8db27bd11ccb1e924e79
size 5751
