version https://git-lfs.github.com/spec/v1
oid sha256:88758b4c88c5c70f5ebe21254dcfef7a6ad093506f6243d03508ba41b237d1c4
size 7034
