version https://git-lfs.github.com/spec/v1
oid sha256:4b575686c502f1b4d0cdbbc50139ed559bc25a0359dd25a880b74d1bda593348
size 4178
